`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/13/2025 01:25:02 AM
// Design Name: 
// Module Name: Imm_gen
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Imm_gen(
    input [31:0] instr,
    output reg [31:0] imm
    );
//wire [6:0] opcode = instr[6:0];
always@(*)
begin
    case(instr[6:0])
    7'b0010011,7'b0000011,7'b1100111 : imm= {{20{instr[31]}},instr[31:20]}; //I-Type JALR type
    7'b0100011: imm={{20{instr[31]}},instr[31:25],instr[11:7]}; //S-Type
    7'b1100011: imm = {{19{instr[31]}}, instr[31], instr[7], instr[30:25], instr[11:8], 1'b0}; // B-type
   // 7'b1101111: imm = {{12{instr[31]}},instr[31:12]}; //JAL-type
    7'b1101111: imm = {{11{instr[31]}}, instr[31], instr[19:12], instr[20], instr[30:21], 1'b0}; // JAL-type
    default: imm = 32'b0;
    endcase
    
   // $display("imm value = %0d", imm);
end
endmodule
